// arm.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module arm (
		output wire [7:0]  buff_export,               //               buff.export
		output wire [7:0]  card_select_export,        //        card_select.export
		input  wire        clk_clk,                   //                clk.clk
		output wire [7:0]  ending_info_export,        //        ending_info.export
		output wire [7:0]  enemy_card_used_export,    //    enemy_card_used.export
		output wire [7:0]  enemy_card_visible_export, // enemy_card_visible.export
		output wire [7:0]  enemy_hp_export,           //           enemy_hp.export
		output wire [7:0]  enemy_shield_export,       //       enemy_shield.export
		output wire [7:0]  initial_screen_export,     //     initial_screen.export
		input  wire [31:0] keycode_export,            //            keycode.export
		output wire [31:0] keycode_reset_export,      //      keycode_reset.export
		output wire [14:0] memory_mem_a,              //             memory.mem_a
		output wire [2:0]  memory_mem_ba,             //                   .mem_ba
		output wire        memory_mem_ck,             //                   .mem_ck
		output wire        memory_mem_ck_n,           //                   .mem_ck_n
		output wire        memory_mem_cke,            //                   .mem_cke
		output wire        memory_mem_cs_n,           //                   .mem_cs_n
		output wire        memory_mem_ras_n,          //                   .mem_ras_n
		output wire        memory_mem_cas_n,          //                   .mem_cas_n
		output wire        memory_mem_we_n,           //                   .mem_we_n
		output wire        memory_mem_reset_n,        //                   .mem_reset_n
		inout  wire [31:0] memory_mem_dq,             //                   .mem_dq
		inout  wire [3:0]  memory_mem_dqs,            //                   .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,          //                   .mem_dqs_n
		output wire        memory_mem_odt,            //                   .mem_odt
		output wire [3:0]  memory_mem_dm,             //                   .mem_dm
		input  wire        memory_oct_rzqin,          //                   .oct_rzqin
		output wire [7:0]  my_card_1_export,          //          my_card_1.export
		output wire [7:0]  my_card_2_export,          //          my_card_2.export
		output wire [7:0]  my_card_3_export,          //          my_card_3.export
		output wire [7:0]  my_card_used_export,       //       my_card_used.export
		output wire [7:0]  my_hp_export,              //              my_hp.export
		output wire [7:0]  my_shield_export,          //          my_shield.export
		input  wire        reset_reset_n,             //              reset.reset_n
		output wire [7:0]  round_export,              //              round.export
		output wire [7:0]  show_instr_export,         //         show_instr.export
		output wire [7:0]  time_export,               //               time.export
		output wire [7:0]  ult_info_export            //           ult_info.export
	);

	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;        // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;          // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;          // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;         // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;            // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;         // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;          // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;            // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;        // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;         // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;         // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;         // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;         // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;          // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;        // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;        // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;           // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;         // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;         // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;         // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;          // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;        // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;          // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;        // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;        // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;         // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;         // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;          // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;          // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;          // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;           // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;            // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;         // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;         // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;        // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;         // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire         mm_interconnect_0_pio_0_s1_chipselect;  // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;    // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;     // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;       // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;   // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire  [31:0] mm_interconnect_0_pio_1_s1_readdata;    // pio_1:readdata -> mm_interconnect_0:pio_1_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_1_s1_address;     // mm_interconnect_0:pio_1_s1_address -> pio_1:address
	wire         mm_interconnect_0_pio_2_s1_chipselect;  // mm_interconnect_0:pio_2_s1_chipselect -> pio_2:chipselect
	wire  [31:0] mm_interconnect_0_pio_2_s1_readdata;    // pio_2:readdata -> mm_interconnect_0:pio_2_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_2_s1_address;     // mm_interconnect_0:pio_2_s1_address -> pio_2:address
	wire         mm_interconnect_0_pio_2_s1_write;       // mm_interconnect_0:pio_2_s1_write -> pio_2:write_n
	wire  [31:0] mm_interconnect_0_pio_2_s1_writedata;   // mm_interconnect_0:pio_2_s1_writedata -> pio_2:writedata
	wire         mm_interconnect_0_pio_3_s1_chipselect;  // mm_interconnect_0:pio_3_s1_chipselect -> pio_3:chipselect
	wire  [31:0] mm_interconnect_0_pio_3_s1_readdata;    // pio_3:readdata -> mm_interconnect_0:pio_3_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_3_s1_address;     // mm_interconnect_0:pio_3_s1_address -> pio_3:address
	wire         mm_interconnect_0_pio_3_s1_write;       // mm_interconnect_0:pio_3_s1_write -> pio_3:write_n
	wire  [31:0] mm_interconnect_0_pio_3_s1_writedata;   // mm_interconnect_0:pio_3_s1_writedata -> pio_3:writedata
	wire         mm_interconnect_0_pio_4_s1_chipselect;  // mm_interconnect_0:pio_4_s1_chipselect -> pio_4:chipselect
	wire  [31:0] mm_interconnect_0_pio_4_s1_readdata;    // pio_4:readdata -> mm_interconnect_0:pio_4_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_4_s1_address;     // mm_interconnect_0:pio_4_s1_address -> pio_4:address
	wire         mm_interconnect_0_pio_4_s1_write;       // mm_interconnect_0:pio_4_s1_write -> pio_4:write_n
	wire  [31:0] mm_interconnect_0_pio_4_s1_writedata;   // mm_interconnect_0:pio_4_s1_writedata -> pio_4:writedata
	wire         mm_interconnect_0_pio_5_s1_chipselect;  // mm_interconnect_0:pio_5_s1_chipselect -> pio_5:chipselect
	wire  [31:0] mm_interconnect_0_pio_5_s1_readdata;    // pio_5:readdata -> mm_interconnect_0:pio_5_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_5_s1_address;     // mm_interconnect_0:pio_5_s1_address -> pio_5:address
	wire         mm_interconnect_0_pio_5_s1_write;       // mm_interconnect_0:pio_5_s1_write -> pio_5:write_n
	wire  [31:0] mm_interconnect_0_pio_5_s1_writedata;   // mm_interconnect_0:pio_5_s1_writedata -> pio_5:writedata
	wire         mm_interconnect_0_pio_6_s1_chipselect;  // mm_interconnect_0:pio_6_s1_chipselect -> pio_6:chipselect
	wire  [31:0] mm_interconnect_0_pio_6_s1_readdata;    // pio_6:readdata -> mm_interconnect_0:pio_6_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_6_s1_address;     // mm_interconnect_0:pio_6_s1_address -> pio_6:address
	wire         mm_interconnect_0_pio_6_s1_write;       // mm_interconnect_0:pio_6_s1_write -> pio_6:write_n
	wire  [31:0] mm_interconnect_0_pio_6_s1_writedata;   // mm_interconnect_0:pio_6_s1_writedata -> pio_6:writedata
	wire         mm_interconnect_0_pio_7_s1_chipselect;  // mm_interconnect_0:pio_7_s1_chipselect -> pio_7:chipselect
	wire  [31:0] mm_interconnect_0_pio_7_s1_readdata;    // pio_7:readdata -> mm_interconnect_0:pio_7_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_7_s1_address;     // mm_interconnect_0:pio_7_s1_address -> pio_7:address
	wire         mm_interconnect_0_pio_7_s1_write;       // mm_interconnect_0:pio_7_s1_write -> pio_7:write_n
	wire  [31:0] mm_interconnect_0_pio_7_s1_writedata;   // mm_interconnect_0:pio_7_s1_writedata -> pio_7:writedata
	wire         mm_interconnect_0_pio_8_s1_chipselect;  // mm_interconnect_0:pio_8_s1_chipselect -> pio_8:chipselect
	wire  [31:0] mm_interconnect_0_pio_8_s1_readdata;    // pio_8:readdata -> mm_interconnect_0:pio_8_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_8_s1_address;     // mm_interconnect_0:pio_8_s1_address -> pio_8:address
	wire         mm_interconnect_0_pio_8_s1_write;       // mm_interconnect_0:pio_8_s1_write -> pio_8:write_n
	wire  [31:0] mm_interconnect_0_pio_8_s1_writedata;   // mm_interconnect_0:pio_8_s1_writedata -> pio_8:writedata
	wire         mm_interconnect_0_pio_9_s1_chipselect;  // mm_interconnect_0:pio_9_s1_chipselect -> pio_9:chipselect
	wire  [31:0] mm_interconnect_0_pio_9_s1_readdata;    // pio_9:readdata -> mm_interconnect_0:pio_9_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_9_s1_address;     // mm_interconnect_0:pio_9_s1_address -> pio_9:address
	wire         mm_interconnect_0_pio_9_s1_write;       // mm_interconnect_0:pio_9_s1_write -> pio_9:write_n
	wire  [31:0] mm_interconnect_0_pio_9_s1_writedata;   // mm_interconnect_0:pio_9_s1_writedata -> pio_9:writedata
	wire         mm_interconnect_0_pio_10_s1_chipselect; // mm_interconnect_0:pio_10_s1_chipselect -> pio_10:chipselect
	wire  [31:0] mm_interconnect_0_pio_10_s1_readdata;   // pio_10:readdata -> mm_interconnect_0:pio_10_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_10_s1_address;    // mm_interconnect_0:pio_10_s1_address -> pio_10:address
	wire         mm_interconnect_0_pio_10_s1_write;      // mm_interconnect_0:pio_10_s1_write -> pio_10:write_n
	wire  [31:0] mm_interconnect_0_pio_10_s1_writedata;  // mm_interconnect_0:pio_10_s1_writedata -> pio_10:writedata
	wire         mm_interconnect_0_pio_11_s1_chipselect; // mm_interconnect_0:pio_11_s1_chipselect -> pio_11:chipselect
	wire  [31:0] mm_interconnect_0_pio_11_s1_readdata;   // pio_11:readdata -> mm_interconnect_0:pio_11_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_11_s1_address;    // mm_interconnect_0:pio_11_s1_address -> pio_11:address
	wire         mm_interconnect_0_pio_11_s1_write;      // mm_interconnect_0:pio_11_s1_write -> pio_11:write_n
	wire  [31:0] mm_interconnect_0_pio_11_s1_writedata;  // mm_interconnect_0:pio_11_s1_writedata -> pio_11:writedata
	wire         mm_interconnect_0_pio_12_s1_chipselect; // mm_interconnect_0:pio_12_s1_chipselect -> pio_12:chipselect
	wire  [31:0] mm_interconnect_0_pio_12_s1_readdata;   // pio_12:readdata -> mm_interconnect_0:pio_12_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_12_s1_address;    // mm_interconnect_0:pio_12_s1_address -> pio_12:address
	wire         mm_interconnect_0_pio_12_s1_write;      // mm_interconnect_0:pio_12_s1_write -> pio_12:write_n
	wire  [31:0] mm_interconnect_0_pio_12_s1_writedata;  // mm_interconnect_0:pio_12_s1_writedata -> pio_12:writedata
	wire         mm_interconnect_0_pio_13_s1_chipselect; // mm_interconnect_0:pio_13_s1_chipselect -> pio_13:chipselect
	wire  [31:0] mm_interconnect_0_pio_13_s1_readdata;   // pio_13:readdata -> mm_interconnect_0:pio_13_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_13_s1_address;    // mm_interconnect_0:pio_13_s1_address -> pio_13:address
	wire         mm_interconnect_0_pio_13_s1_write;      // mm_interconnect_0:pio_13_s1_write -> pio_13:write_n
	wire  [31:0] mm_interconnect_0_pio_13_s1_writedata;  // mm_interconnect_0:pio_13_s1_writedata -> pio_13:writedata
	wire         mm_interconnect_0_pio_14_s1_chipselect; // mm_interconnect_0:pio_14_s1_chipselect -> pio_14:chipselect
	wire  [31:0] mm_interconnect_0_pio_14_s1_readdata;   // pio_14:readdata -> mm_interconnect_0:pio_14_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_14_s1_address;    // mm_interconnect_0:pio_14_s1_address -> pio_14:address
	wire         mm_interconnect_0_pio_14_s1_write;      // mm_interconnect_0:pio_14_s1_write -> pio_14:write_n
	wire  [31:0] mm_interconnect_0_pio_14_s1_writedata;  // mm_interconnect_0:pio_14_s1_writedata -> pio_14:writedata
	wire         mm_interconnect_0_pio_15_s1_chipselect; // mm_interconnect_0:pio_15_s1_chipselect -> pio_15:chipselect
	wire  [31:0] mm_interconnect_0_pio_15_s1_readdata;   // pio_15:readdata -> mm_interconnect_0:pio_15_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_15_s1_address;    // mm_interconnect_0:pio_15_s1_address -> pio_15:address
	wire         mm_interconnect_0_pio_15_s1_write;      // mm_interconnect_0:pio_15_s1_write -> pio_15:write_n
	wire  [31:0] mm_interconnect_0_pio_15_s1_writedata;  // mm_interconnect_0:pio_15_s1_writedata -> pio_15:writedata
	wire         mm_interconnect_0_pio_16_s1_chipselect; // mm_interconnect_0:pio_16_s1_chipselect -> pio_16:chipselect
	wire  [31:0] mm_interconnect_0_pio_16_s1_readdata;   // pio_16:readdata -> mm_interconnect_0:pio_16_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_16_s1_address;    // mm_interconnect_0:pio_16_s1_address -> pio_16:address
	wire         mm_interconnect_0_pio_16_s1_write;      // mm_interconnect_0:pio_16_s1_write -> pio_16:write_n
	wire  [31:0] mm_interconnect_0_pio_16_s1_writedata;  // mm_interconnect_0:pio_16_s1_writedata -> pio_16:writedata
	wire         mm_interconnect_0_pio_17_s1_chipselect; // mm_interconnect_0:pio_17_s1_chipselect -> pio_17:chipselect
	wire  [31:0] mm_interconnect_0_pio_17_s1_readdata;   // pio_17:readdata -> mm_interconnect_0:pio_17_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_17_s1_address;    // mm_interconnect_0:pio_17_s1_address -> pio_17:address
	wire         mm_interconnect_0_pio_17_s1_write;      // mm_interconnect_0:pio_17_s1_write -> pio_17:write_n
	wire  [31:0] mm_interconnect_0_pio_17_s1_writedata;  // mm_interconnect_0:pio_17_s1_writedata -> pio_17:writedata
	wire         mm_interconnect_0_pio_18_s1_chipselect; // mm_interconnect_0:pio_18_s1_chipselect -> pio_18:chipselect
	wire  [31:0] mm_interconnect_0_pio_18_s1_readdata;   // pio_18:readdata -> mm_interconnect_0:pio_18_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_18_s1_address;    // mm_interconnect_0:pio_18_s1_address -> pio_18:address
	wire         mm_interconnect_0_pio_18_s1_write;      // mm_interconnect_0:pio_18_s1_write -> pio_18:write_n
	wire  [31:0] mm_interconnect_0_pio_18_s1_writedata;  // mm_interconnect_0:pio_18_s1_writedata -> pio_18:writedata
	wire         mm_interconnect_0_pio_19_s1_chipselect; // mm_interconnect_0:pio_19_s1_chipselect -> pio_19:chipselect
	wire  [31:0] mm_interconnect_0_pio_19_s1_readdata;   // pio_19:readdata -> mm_interconnect_0:pio_19_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_19_s1_address;    // mm_interconnect_0:pio_19_s1_address -> pio_19:address
	wire         mm_interconnect_0_pio_19_s1_write;      // mm_interconnect_0:pio_19_s1_write -> pio_19:write_n
	wire  [31:0] mm_interconnect_0_pio_19_s1_writedata;  // mm_interconnect_0:pio_19_s1_writedata -> pio_19:writedata
	wire         rst_controller_reset_out_reset;         // rst_controller:reset_out -> [mm_interconnect_0:pio_0_reset_reset_bridge_in_reset_reset, pio_0:reset_n, pio_10:reset_n, pio_11:reset_n, pio_12:reset_n, pio_13:reset_n, pio_14:reset_n, pio_15:reset_n, pio_16:reset_n, pio_17:reset_n, pio_18:reset_n, pio_19:reset_n, pio_1:reset_n, pio_2:reset_n, pio_3:reset_n, pio_4:reset_n, pio_5:reset_n, pio_6:reset_n, pio_7:reset_n, pio_8:reset_n, pio_9:reset_n]
	wire         rst_controller_001_reset_out_reset;     // rst_controller_001:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         hps_0_h2f_reset_reset;                  // hps_0:h2f_rst_n -> rst_controller_001:reset_in0

	arm_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (3)
	) hps_0 (
		.mem_a          (memory_mem_a),                    //            memory.mem_a
		.mem_ba         (memory_mem_ba),                   //                  .mem_ba
		.mem_ck         (memory_mem_ck),                   //                  .mem_ck
		.mem_ck_n       (memory_mem_ck_n),                 //                  .mem_ck_n
		.mem_cke        (memory_mem_cke),                  //                  .mem_cke
		.mem_cs_n       (memory_mem_cs_n),                 //                  .mem_cs_n
		.mem_ras_n      (memory_mem_ras_n),                //                  .mem_ras_n
		.mem_cas_n      (memory_mem_cas_n),                //                  .mem_cas_n
		.mem_we_n       (memory_mem_we_n),                 //                  .mem_we_n
		.mem_reset_n    (memory_mem_reset_n),              //                  .mem_reset_n
		.mem_dq         (memory_mem_dq),                   //                  .mem_dq
		.mem_dqs        (memory_mem_dqs),                  //                  .mem_dqs
		.mem_dqs_n      (memory_mem_dqs_n),                //                  .mem_dqs_n
		.mem_odt        (memory_mem_odt),                  //                  .mem_odt
		.mem_dm         (memory_mem_dm),                   //                  .mem_dm
		.oct_rzqin      (memory_oct_rzqin),                //                  .oct_rzqin
		.h2f_rst_n      (hps_0_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_axi_clk    (clk_clk),                         //     h2f_axi_clock.clk
		.h2f_AWID       (),                                //    h2f_axi_master.awid
		.h2f_AWADDR     (),                                //                  .awaddr
		.h2f_AWLEN      (),                                //                  .awlen
		.h2f_AWSIZE     (),                                //                  .awsize
		.h2f_AWBURST    (),                                //                  .awburst
		.h2f_AWLOCK     (),                                //                  .awlock
		.h2f_AWCACHE    (),                                //                  .awcache
		.h2f_AWPROT     (),                                //                  .awprot
		.h2f_AWVALID    (),                                //                  .awvalid
		.h2f_AWREADY    (),                                //                  .awready
		.h2f_WID        (),                                //                  .wid
		.h2f_WDATA      (),                                //                  .wdata
		.h2f_WSTRB      (),                                //                  .wstrb
		.h2f_WLAST      (),                                //                  .wlast
		.h2f_WVALID     (),                                //                  .wvalid
		.h2f_WREADY     (),                                //                  .wready
		.h2f_BID        (),                                //                  .bid
		.h2f_BRESP      (),                                //                  .bresp
		.h2f_BVALID     (),                                //                  .bvalid
		.h2f_BREADY     (),                                //                  .bready
		.h2f_ARID       (),                                //                  .arid
		.h2f_ARADDR     (),                                //                  .araddr
		.h2f_ARLEN      (),                                //                  .arlen
		.h2f_ARSIZE     (),                                //                  .arsize
		.h2f_ARBURST    (),                                //                  .arburst
		.h2f_ARLOCK     (),                                //                  .arlock
		.h2f_ARCACHE    (),                                //                  .arcache
		.h2f_ARPROT     (),                                //                  .arprot
		.h2f_ARVALID    (),                                //                  .arvalid
		.h2f_ARREADY    (),                                //                  .arready
		.h2f_RID        (),                                //                  .rid
		.h2f_RDATA      (),                                //                  .rdata
		.h2f_RRESP      (),                                //                  .rresp
		.h2f_RLAST      (),                                //                  .rlast
		.h2f_RVALID     (),                                //                  .rvalid
		.h2f_RREADY     (),                                //                  .rready
		.f2h_axi_clk    (clk_clk),                         //     f2h_axi_clock.clk
		.f2h_AWID       (),                                //     f2h_axi_slave.awid
		.f2h_AWADDR     (),                                //                  .awaddr
		.f2h_AWLEN      (),                                //                  .awlen
		.f2h_AWSIZE     (),                                //                  .awsize
		.f2h_AWBURST    (),                                //                  .awburst
		.f2h_AWLOCK     (),                                //                  .awlock
		.f2h_AWCACHE    (),                                //                  .awcache
		.f2h_AWPROT     (),                                //                  .awprot
		.f2h_AWVALID    (),                                //                  .awvalid
		.f2h_AWREADY    (),                                //                  .awready
		.f2h_AWUSER     (),                                //                  .awuser
		.f2h_WID        (),                                //                  .wid
		.f2h_WDATA      (),                                //                  .wdata
		.f2h_WSTRB      (),                                //                  .wstrb
		.f2h_WLAST      (),                                //                  .wlast
		.f2h_WVALID     (),                                //                  .wvalid
		.f2h_WREADY     (),                                //                  .wready
		.f2h_BID        (),                                //                  .bid
		.f2h_BRESP      (),                                //                  .bresp
		.f2h_BVALID     (),                                //                  .bvalid
		.f2h_BREADY     (),                                //                  .bready
		.f2h_ARID       (),                                //                  .arid
		.f2h_ARADDR     (),                                //                  .araddr
		.f2h_ARLEN      (),                                //                  .arlen
		.f2h_ARSIZE     (),                                //                  .arsize
		.f2h_ARBURST    (),                                //                  .arburst
		.f2h_ARLOCK     (),                                //                  .arlock
		.f2h_ARCACHE    (),                                //                  .arcache
		.f2h_ARPROT     (),                                //                  .arprot
		.f2h_ARVALID    (),                                //                  .arvalid
		.f2h_ARREADY    (),                                //                  .arready
		.f2h_ARUSER     (),                                //                  .aruser
		.f2h_RID        (),                                //                  .rid
		.f2h_RDATA      (),                                //                  .rdata
		.f2h_RRESP      (),                                //                  .rresp
		.f2h_RLAST      (),                                //                  .rlast
		.f2h_RVALID     (),                                //                  .rvalid
		.f2h_RREADY     (),                                //                  .rready
		.h2f_lw_axi_clk (clk_clk),                         //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID    (hps_0_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR  (hps_0_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN   (hps_0_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE  (hps_0_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST (hps_0_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK  (hps_0_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE (hps_0_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT  (hps_0_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID (hps_0_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY (hps_0_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID     (hps_0_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA   (hps_0_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB   (hps_0_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST   (hps_0_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID  (hps_0_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY  (hps_0_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID     (hps_0_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP   (hps_0_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID  (hps_0_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY  (hps_0_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID    (hps_0_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR  (hps_0_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN   (hps_0_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE  (hps_0_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST (hps_0_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK  (hps_0_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE (hps_0_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT  (hps_0_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID (hps_0_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY (hps_0_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID     (hps_0_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA   (hps_0_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP   (hps_0_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST   (hps_0_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID  (hps_0_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY  (hps_0_h2f_lw_axi_master_rready)   //                  .rready
	);

	arm_pio_0 pio_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (initial_screen_export)                  // external_connection.export
	);

	arm_pio_1 pio_1 (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_pio_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_1_s1_readdata), //                    .readdata
		.in_port  (keycode_export)                       // external_connection.export
	);

	arm_pio_0 pio_10 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_pio_10_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_10_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_10_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_10_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_10_s1_readdata),   //                    .readdata
		.out_port   (my_hp_export)                            // external_connection.export
	);

	arm_pio_0 pio_11 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_pio_11_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_11_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_11_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_11_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_11_s1_readdata),   //                    .readdata
		.out_port   (my_shield_export)                        // external_connection.export
	);

	arm_pio_0 pio_12 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_pio_12_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_12_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_12_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_12_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_12_s1_readdata),   //                    .readdata
		.out_port   (time_export)                             // external_connection.export
	);

	arm_pio_0 pio_13 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_pio_13_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_13_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_13_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_13_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_13_s1_readdata),   //                    .readdata
		.out_port   (round_export)                            // external_connection.export
	);

	arm_pio_0 pio_14 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_pio_14_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_14_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_14_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_14_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_14_s1_readdata),   //                    .readdata
		.out_port   (enemy_hp_export)                         // external_connection.export
	);

	arm_pio_0 pio_15 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_pio_15_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_15_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_15_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_15_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_15_s1_readdata),   //                    .readdata
		.out_port   (enemy_shield_export)                     // external_connection.export
	);

	arm_pio_0 pio_16 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_pio_16_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_16_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_16_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_16_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_16_s1_readdata),   //                    .readdata
		.out_port   (buff_export)                             // external_connection.export
	);

	arm_pio_0 pio_17 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_pio_17_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_17_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_17_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_17_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_17_s1_readdata),   //                    .readdata
		.out_port   (ult_info_export)                         // external_connection.export
	);

	arm_pio_0 pio_18 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_pio_18_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_18_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_18_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_18_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_18_s1_readdata),   //                    .readdata
		.out_port   (ending_info_export)                      // external_connection.export
	);

	arm_pio_0 pio_19 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_pio_19_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_19_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_19_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_19_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_19_s1_readdata),   //                    .readdata
		.out_port   (show_instr_export)                       // external_connection.export
	);

	arm_pio_2 pio_2 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_2_s1_readdata),   //                    .readdata
		.out_port   (keycode_reset_export)                   // external_connection.export
	);

	arm_pio_0 pio_3 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_3_s1_readdata),   //                    .readdata
		.out_port   (card_select_export)                     // external_connection.export
	);

	arm_pio_0 pio_4 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_4_s1_readdata),   //                    .readdata
		.out_port   (my_card_1_export)                       // external_connection.export
	);

	arm_pio_0 pio_5 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_5_s1_readdata),   //                    .readdata
		.out_port   (my_card_2_export)                       // external_connection.export
	);

	arm_pio_0 pio_6 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_6_s1_readdata),   //                    .readdata
		.out_port   (my_card_3_export)                       // external_connection.export
	);

	arm_pio_0 pio_7 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_7_s1_readdata),   //                    .readdata
		.out_port   (my_card_used_export)                    // external_connection.export
	);

	arm_pio_0 pio_8 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_8_s1_readdata),   //                    .readdata
		.out_port   (enemy_card_used_export)                 // external_connection.export
	);

	arm_pio_0 pio_9 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_9_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_9_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_9_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_9_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_9_s1_readdata),   //                    .readdata
		.out_port   (enemy_card_visible_export)              // external_connection.export
	);

	arm_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),           //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),         //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),          //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),         //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),        //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),         //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),        //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),         //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),        //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),        //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),            //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),          //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),          //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),          //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),         //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),         //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),            //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),          //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),         //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),         //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),           //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),         //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),          //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),         //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),        //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),         //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),        //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),         //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),        //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),        //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),            //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),          //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),          //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),          //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),         //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),         //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                //                                                     clk_0_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),     // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.pio_0_reset_reset_bridge_in_reset_reset                             (rst_controller_reset_out_reset),         //                             pio_0_reset_reset_bridge_in_reset.reset
		.pio_0_s1_address                                                    (mm_interconnect_0_pio_0_s1_address),     //                                                      pio_0_s1.address
		.pio_0_s1_write                                                      (mm_interconnect_0_pio_0_s1_write),       //                                                              .write
		.pio_0_s1_readdata                                                   (mm_interconnect_0_pio_0_s1_readdata),    //                                                              .readdata
		.pio_0_s1_writedata                                                  (mm_interconnect_0_pio_0_s1_writedata),   //                                                              .writedata
		.pio_0_s1_chipselect                                                 (mm_interconnect_0_pio_0_s1_chipselect),  //                                                              .chipselect
		.pio_1_s1_address                                                    (mm_interconnect_0_pio_1_s1_address),     //                                                      pio_1_s1.address
		.pio_1_s1_readdata                                                   (mm_interconnect_0_pio_1_s1_readdata),    //                                                              .readdata
		.pio_10_s1_address                                                   (mm_interconnect_0_pio_10_s1_address),    //                                                     pio_10_s1.address
		.pio_10_s1_write                                                     (mm_interconnect_0_pio_10_s1_write),      //                                                              .write
		.pio_10_s1_readdata                                                  (mm_interconnect_0_pio_10_s1_readdata),   //                                                              .readdata
		.pio_10_s1_writedata                                                 (mm_interconnect_0_pio_10_s1_writedata),  //                                                              .writedata
		.pio_10_s1_chipselect                                                (mm_interconnect_0_pio_10_s1_chipselect), //                                                              .chipselect
		.pio_11_s1_address                                                   (mm_interconnect_0_pio_11_s1_address),    //                                                     pio_11_s1.address
		.pio_11_s1_write                                                     (mm_interconnect_0_pio_11_s1_write),      //                                                              .write
		.pio_11_s1_readdata                                                  (mm_interconnect_0_pio_11_s1_readdata),   //                                                              .readdata
		.pio_11_s1_writedata                                                 (mm_interconnect_0_pio_11_s1_writedata),  //                                                              .writedata
		.pio_11_s1_chipselect                                                (mm_interconnect_0_pio_11_s1_chipselect), //                                                              .chipselect
		.pio_12_s1_address                                                   (mm_interconnect_0_pio_12_s1_address),    //                                                     pio_12_s1.address
		.pio_12_s1_write                                                     (mm_interconnect_0_pio_12_s1_write),      //                                                              .write
		.pio_12_s1_readdata                                                  (mm_interconnect_0_pio_12_s1_readdata),   //                                                              .readdata
		.pio_12_s1_writedata                                                 (mm_interconnect_0_pio_12_s1_writedata),  //                                                              .writedata
		.pio_12_s1_chipselect                                                (mm_interconnect_0_pio_12_s1_chipselect), //                                                              .chipselect
		.pio_13_s1_address                                                   (mm_interconnect_0_pio_13_s1_address),    //                                                     pio_13_s1.address
		.pio_13_s1_write                                                     (mm_interconnect_0_pio_13_s1_write),      //                                                              .write
		.pio_13_s1_readdata                                                  (mm_interconnect_0_pio_13_s1_readdata),   //                                                              .readdata
		.pio_13_s1_writedata                                                 (mm_interconnect_0_pio_13_s1_writedata),  //                                                              .writedata
		.pio_13_s1_chipselect                                                (mm_interconnect_0_pio_13_s1_chipselect), //                                                              .chipselect
		.pio_14_s1_address                                                   (mm_interconnect_0_pio_14_s1_address),    //                                                     pio_14_s1.address
		.pio_14_s1_write                                                     (mm_interconnect_0_pio_14_s1_write),      //                                                              .write
		.pio_14_s1_readdata                                                  (mm_interconnect_0_pio_14_s1_readdata),   //                                                              .readdata
		.pio_14_s1_writedata                                                 (mm_interconnect_0_pio_14_s1_writedata),  //                                                              .writedata
		.pio_14_s1_chipselect                                                (mm_interconnect_0_pio_14_s1_chipselect), //                                                              .chipselect
		.pio_15_s1_address                                                   (mm_interconnect_0_pio_15_s1_address),    //                                                     pio_15_s1.address
		.pio_15_s1_write                                                     (mm_interconnect_0_pio_15_s1_write),      //                                                              .write
		.pio_15_s1_readdata                                                  (mm_interconnect_0_pio_15_s1_readdata),   //                                                              .readdata
		.pio_15_s1_writedata                                                 (mm_interconnect_0_pio_15_s1_writedata),  //                                                              .writedata
		.pio_15_s1_chipselect                                                (mm_interconnect_0_pio_15_s1_chipselect), //                                                              .chipselect
		.pio_16_s1_address                                                   (mm_interconnect_0_pio_16_s1_address),    //                                                     pio_16_s1.address
		.pio_16_s1_write                                                     (mm_interconnect_0_pio_16_s1_write),      //                                                              .write
		.pio_16_s1_readdata                                                  (mm_interconnect_0_pio_16_s1_readdata),   //                                                              .readdata
		.pio_16_s1_writedata                                                 (mm_interconnect_0_pio_16_s1_writedata),  //                                                              .writedata
		.pio_16_s1_chipselect                                                (mm_interconnect_0_pio_16_s1_chipselect), //                                                              .chipselect
		.pio_17_s1_address                                                   (mm_interconnect_0_pio_17_s1_address),    //                                                     pio_17_s1.address
		.pio_17_s1_write                                                     (mm_interconnect_0_pio_17_s1_write),      //                                                              .write
		.pio_17_s1_readdata                                                  (mm_interconnect_0_pio_17_s1_readdata),   //                                                              .readdata
		.pio_17_s1_writedata                                                 (mm_interconnect_0_pio_17_s1_writedata),  //                                                              .writedata
		.pio_17_s1_chipselect                                                (mm_interconnect_0_pio_17_s1_chipselect), //                                                              .chipselect
		.pio_18_s1_address                                                   (mm_interconnect_0_pio_18_s1_address),    //                                                     pio_18_s1.address
		.pio_18_s1_write                                                     (mm_interconnect_0_pio_18_s1_write),      //                                                              .write
		.pio_18_s1_readdata                                                  (mm_interconnect_0_pio_18_s1_readdata),   //                                                              .readdata
		.pio_18_s1_writedata                                                 (mm_interconnect_0_pio_18_s1_writedata),  //                                                              .writedata
		.pio_18_s1_chipselect                                                (mm_interconnect_0_pio_18_s1_chipselect), //                                                              .chipselect
		.pio_19_s1_address                                                   (mm_interconnect_0_pio_19_s1_address),    //                                                     pio_19_s1.address
		.pio_19_s1_write                                                     (mm_interconnect_0_pio_19_s1_write),      //                                                              .write
		.pio_19_s1_readdata                                                  (mm_interconnect_0_pio_19_s1_readdata),   //                                                              .readdata
		.pio_19_s1_writedata                                                 (mm_interconnect_0_pio_19_s1_writedata),  //                                                              .writedata
		.pio_19_s1_chipselect                                                (mm_interconnect_0_pio_19_s1_chipselect), //                                                              .chipselect
		.pio_2_s1_address                                                    (mm_interconnect_0_pio_2_s1_address),     //                                                      pio_2_s1.address
		.pio_2_s1_write                                                      (mm_interconnect_0_pio_2_s1_write),       //                                                              .write
		.pio_2_s1_readdata                                                   (mm_interconnect_0_pio_2_s1_readdata),    //                                                              .readdata
		.pio_2_s1_writedata                                                  (mm_interconnect_0_pio_2_s1_writedata),   //                                                              .writedata
		.pio_2_s1_chipselect                                                 (mm_interconnect_0_pio_2_s1_chipselect),  //                                                              .chipselect
		.pio_3_s1_address                                                    (mm_interconnect_0_pio_3_s1_address),     //                                                      pio_3_s1.address
		.pio_3_s1_write                                                      (mm_interconnect_0_pio_3_s1_write),       //                                                              .write
		.pio_3_s1_readdata                                                   (mm_interconnect_0_pio_3_s1_readdata),    //                                                              .readdata
		.pio_3_s1_writedata                                                  (mm_interconnect_0_pio_3_s1_writedata),   //                                                              .writedata
		.pio_3_s1_chipselect                                                 (mm_interconnect_0_pio_3_s1_chipselect),  //                                                              .chipselect
		.pio_4_s1_address                                                    (mm_interconnect_0_pio_4_s1_address),     //                                                      pio_4_s1.address
		.pio_4_s1_write                                                      (mm_interconnect_0_pio_4_s1_write),       //                                                              .write
		.pio_4_s1_readdata                                                   (mm_interconnect_0_pio_4_s1_readdata),    //                                                              .readdata
		.pio_4_s1_writedata                                                  (mm_interconnect_0_pio_4_s1_writedata),   //                                                              .writedata
		.pio_4_s1_chipselect                                                 (mm_interconnect_0_pio_4_s1_chipselect),  //                                                              .chipselect
		.pio_5_s1_address                                                    (mm_interconnect_0_pio_5_s1_address),     //                                                      pio_5_s1.address
		.pio_5_s1_write                                                      (mm_interconnect_0_pio_5_s1_write),       //                                                              .write
		.pio_5_s1_readdata                                                   (mm_interconnect_0_pio_5_s1_readdata),    //                                                              .readdata
		.pio_5_s1_writedata                                                  (mm_interconnect_0_pio_5_s1_writedata),   //                                                              .writedata
		.pio_5_s1_chipselect                                                 (mm_interconnect_0_pio_5_s1_chipselect),  //                                                              .chipselect
		.pio_6_s1_address                                                    (mm_interconnect_0_pio_6_s1_address),     //                                                      pio_6_s1.address
		.pio_6_s1_write                                                      (mm_interconnect_0_pio_6_s1_write),       //                                                              .write
		.pio_6_s1_readdata                                                   (mm_interconnect_0_pio_6_s1_readdata),    //                                                              .readdata
		.pio_6_s1_writedata                                                  (mm_interconnect_0_pio_6_s1_writedata),   //                                                              .writedata
		.pio_6_s1_chipselect                                                 (mm_interconnect_0_pio_6_s1_chipselect),  //                                                              .chipselect
		.pio_7_s1_address                                                    (mm_interconnect_0_pio_7_s1_address),     //                                                      pio_7_s1.address
		.pio_7_s1_write                                                      (mm_interconnect_0_pio_7_s1_write),       //                                                              .write
		.pio_7_s1_readdata                                                   (mm_interconnect_0_pio_7_s1_readdata),    //                                                              .readdata
		.pio_7_s1_writedata                                                  (mm_interconnect_0_pio_7_s1_writedata),   //                                                              .writedata
		.pio_7_s1_chipselect                                                 (mm_interconnect_0_pio_7_s1_chipselect),  //                                                              .chipselect
		.pio_8_s1_address                                                    (mm_interconnect_0_pio_8_s1_address),     //                                                      pio_8_s1.address
		.pio_8_s1_write                                                      (mm_interconnect_0_pio_8_s1_write),       //                                                              .write
		.pio_8_s1_readdata                                                   (mm_interconnect_0_pio_8_s1_readdata),    //                                                              .readdata
		.pio_8_s1_writedata                                                  (mm_interconnect_0_pio_8_s1_writedata),   //                                                              .writedata
		.pio_8_s1_chipselect                                                 (mm_interconnect_0_pio_8_s1_chipselect),  //                                                              .chipselect
		.pio_9_s1_address                                                    (mm_interconnect_0_pio_9_s1_address),     //                                                      pio_9_s1.address
		.pio_9_s1_write                                                      (mm_interconnect_0_pio_9_s1_write),       //                                                              .write
		.pio_9_s1_readdata                                                   (mm_interconnect_0_pio_9_s1_readdata),    //                                                              .readdata
		.pio_9_s1_writedata                                                  (mm_interconnect_0_pio_9_s1_writedata),   //                                                              .writedata
		.pio_9_s1_chipselect                                                 (mm_interconnect_0_pio_9_s1_chipselect)   //                                                              .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
